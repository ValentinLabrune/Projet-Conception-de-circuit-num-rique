library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity MemInstruction is
    port(
        clock_IN : in std_logic;
        reset_IN : in std_logic;

        SEL_FCT_OUT : out std_logic_vector (3 downto 0);
        SEL_ROUTE_OUT : out std_logic_vector (3 downto 0);
        SEL_OUT_OUT : out std_logic_vector (1 downto 0)
    );
end MemInstruction;

architecture MemInstruction_Arch of MemInstruction is

    -- memoire
    type memory is array (0 to 127) of std_logic_vector (9 downto 0); 
    signal pointeur : integer range 0 to 127 := 0;

    constant MemInstruction : memory := (
        ("0000000000"),  -- pointeur : 0

        -- operation 1
        ("0000011100"), -- pointeur : 1
        ("0000111100"), -- 2
        ("1101000011"), -- 3

        -- operation 2
        ("0000011100"), -- 4
        ("0000111100"), -- 5
        ("1011000000"), -- 6
        ("0000100000"), -- 7
        ("0000011100"), -- 8
        ("0101000000"), -- 9
        ("0000010100"), -- 10
        ("0000100100"), -- 11
        ("1001000011"), -- 12

        -- opération 3

        ("0000011100"), -- 13
        ("0000111100"), -- 14
        ("0111000000"), -- 15
        ("0000100000"), -- 16
        ("0000011100"), -- 17
        ("0000111100"), -- 18
        ("0111000000"), -- 19
        ("0000010100"), -- 20
        ("0000100100"), -- 21
        ("1000000011"), -- 22

        -- remplissage de la memoire de 0
        ("0000000000"), -- 23
        ("0000000000"), -- 24
        ("0000000000"), -- 25
        ("0000000000"), -- 26
        ("0000000000"), -- 27
        ("0000000000"), -- 28
        ("0000000000"), -- 29
        ("0000000000"), -- 30
        ("0000000000"), -- 31
        ("0000000000"), -- 32
        ("0000000000"), -- 33
        ("0000000000"), -- 34
        ("0000000000"), -- 35
        ("0000000000"), -- 36
        ("0000000000"), -- 37
        ("0000000000"), -- 38
        ("0000000000"), -- 39
        ("0000000000"), -- 40
        ("0000000000"), -- 41
        ("0000000000"), -- 42
        ("0000000000"), -- 43
        ("0000000000"), -- 44
        ("0000000000"), -- 45
        ("0000000000"), -- 46
        ("0000000000"), -- 47
        ("0000000000"), -- 48
        ("0000000000"), -- 49
        ("0000000000"), -- 50
        ("0000000000"), -- 51
        ("0000000000"), -- 52
        ("0000000000"), -- 53
        ("0000000000"), -- 54
        ("0000000000"), -- 55
        ("0000000000"), -- 56
        ("0000000000"), -- 57
        ("0000000000"), -- 58
        ("0000000000"), -- 59
        ("0000000000"), -- 60
        ("0000000000"), -- 61
        ("0000000000"), -- 62
        ("0000000000"), -- 63
        ("0000000000"), -- 64
        ("0000000000"), -- 65
        ("0000000000"), -- 66
        ("0000000000"), -- 67
        ("0000000000"), -- 68
        ("0000000000"), -- 69
        ("0000000000"), -- 70
        ("0000000000"), -- 71
        ("0000000000"), -- 72
        ("0000000000"), -- 73
        ("0000000000"), -- 74
        ("0000000000"), -- 75
        ("0000000000"), -- 76
        ("0000000000"), -- 77
        ("0000000000"), -- 78
        ("0000000000"), -- 79
        ("0000000000"), -- 80
        ("0000000000"), -- 81
        ("0000000000"), -- 82
        ("0000000000"), -- 83
        ("0000000000"), -- 84
        ("0000000000"), -- 85
        ("0000000000"), -- 86
        ("0000000000"), -- 87
        ("0000000000"), -- 88
        ("0000000000"), -- 89
        ("0000000000"), -- 90
        ("0000000000"), -- 91
        ("0000000000"), -- 92
        ("0000000000"), -- 93
        ("0000000000"), -- 94
        ("0000000000"), -- 95
        ("0000000000"), -- 96
        ("0000000000"), -- 97
        ("0000000000"), -- 98
        ("0000000000"), -- 99
        ("0000000000"), -- 100
        ("0000000000"), -- 101
        ("0000000000"), -- 102
        ("0000000000"), -- 103
        ("0000000000"), -- 104
        ("0000000000"), -- 105
        ("0000000000"), -- 106
        ("0000000000"), -- 107
        ("0000000000"), -- 108
        ("0000000000"), -- 109
        ("0000000000"), -- 110
        ("0000000000"), -- 111
        ("0000000000"), -- 112
        ("0000000000"), -- 113
        ("0000000000"), -- 114
        ("0000000000"), -- 115
        ("0000000000"), -- 116
        ("0000000000"), -- 117
        ("0000000000"), -- 118
        ("0000000000"), -- 119
        ("0000000000"), -- 120
        ("0000000000"), -- 121
        ("0000000000"), -- 122
        ("0000000000"), -- 123
        ("0000000000"), -- 124
        ("0000000000"), -- 125
        ("0000000000"), -- 126
        ("0000000000") -- 127
        

    );

begin

    process (clock_IN)
    begin
        if (rising_edge(clock_IN)) then
            if (reset_IN = '1') then
                pointeur <= 0;
            else
                pointeur <= pointeur + 1;
            end if;
        end if;
    end process;

    SEL_FCT_OUT <= MemInstruction(pointeur)(9 downto 6);
    SEL_ROUTE_OUT <= MemInstruction(pointeur)(5 downto 2);
    SEL_OUT_OUT <= MemInstruction(pointeur)(1 downto 0);

end MemInstruction_Arch;
    
